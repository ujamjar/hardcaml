module hello_world ();

  initial begin
    $hello;
  end

endmodule

